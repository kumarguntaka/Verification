/**************************************************************************
***                                                                     *** 
***         Kumar Sai Reddy, Fall, 2023									*** 
***                                                                     *** 
*************************************************************************** 
***  Filename: design.sv    Created by Kumar Sai Reddy, 3/29/2023       ***  
***  Version                Version V0p1                                ***  
***  Status                 Tested                                      ***  
***************************************************************************/

package tw_factor_ifft_pkg;

parameter real W128R[0:63]={1.0000000000000000,0.9987954562051724,0.9951847266721969,0.9891765099647810,0.9807852804032304,0.9700312531945440,0.9569403357322088,0.9415440651830208,0.9238795325112867,0.9039892931234433,0.8819212643483550,0.8577286100002721,0.8314696123025452,0.8032075314806449,0.7730104533627370,0.7409511253549591,0.7071067811865476,0.6715589548470183,0.6343932841636455,0.5956993044924335,0.5555702330196023,0.5141027441932217,0.4713967368259978,0.4275550934302822,0.3826834323650898,0.3368898533922201,0.2902846772544623,0.2429801799032640,0.1950903220161283,0.1467304744553617,0.0980171403295608,0.0490676743274181,0.0000000000000001,-0.0490676743274180,-0.0980171403295606,-0.1467304744553616,-0.1950903220161282,-0.2429801799032639,-0.2902846772544622,-0.3368898533922199,-0.3826834323650897,-0.4275550934302819,-0.4713967368259977,-0.5141027441932217,-0.5555702330196020,-0.5956993044924334,-0.6343932841636454,-0.6715589548470184,-0.7071067811865475,-0.7409511253549589,-0.7730104533627370,-0.8032075314806448,-0.8314696123025453,-0.8577286100002720,-0.8819212643483549,-0.9039892931234433,-0.9238795325112867,-0.9415440651830207,-0.9569403357322088,-0.9700312531945440,-0.9807852804032304,-0.9891765099647810,-0.9951847266721968,-0.9987954562051724};
parameter real W128I[0:63]={0.0000000000000000,0.0490676743274180,0.0980171403295606,0.1467304744553617,0.1950903220161282,0.2429801799032639,0.2902846772544623,0.3368898533922201,0.3826834323650898,0.4275550934302821,0.4713967368259976,0.5141027441932217,0.5555702330196022,0.5956993044924334,0.6343932841636455,0.6715589548470183,0.7071067811865475,0.7409511253549591,0.7730104533627370,0.8032075314806448,0.8314696123025452,0.8577286100002721,0.8819212643483549,0.9039892931234433,0.9238795325112867,0.9415440651830208,0.9569403357322089,0.9700312531945440,0.9807852804032304,0.9891765099647810,0.9951847266721968,0.9987954562051724,1.0000000000000000,0.9987954562051724,0.9951847266721969,0.9891765099647810,0.9807852804032304,0.9700312531945440,0.9569403357322089,0.9415440651830208,0.9238795325112867,0.9039892931234434,0.8819212643483550,0.8577286100002721,0.8314696123025455,0.8032075314806449,0.7730104533627371,0.7409511253549590,0.7071067811865476,0.6715589548470186,0.6343932841636455,0.5956993044924335,0.5555702330196022,0.5141027441932218,0.4713967368259979,0.4275550934302820,0.3826834323650899,0.3368898533922203,0.2902846772544624,0.2429801799032641,0.1950903220161286,0.1467304744553618,0.0980171403295608,0.0490676743274180};

endpackage